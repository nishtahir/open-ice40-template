module Top (
    input clk
);

endmodule