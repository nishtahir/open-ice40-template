module Top (
    input clk,
    output LED_G
);

assign LED_G = clk;

endmodule